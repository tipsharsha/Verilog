module parity(

input x,y,z,

output F 
);

xor X (F,x,y,z);  

endmodule